module speed_sel(
		clk,rst_n,


);

input clk;			// 50MHz��ʱ��
input rst_n;		//�͵�ƽ��λ�ź�


/*
parameter bps9600 = 5207;
parameter bps9600_2 = 2603;


*/







endmodule