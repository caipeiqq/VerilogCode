module diplay(
	clk,


);